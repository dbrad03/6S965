module data_framer #
	(
		parameter integer C_M00_AXIS_TDATA_WIDTH	= 32
	)
	(
        input wire pixel_clk,
        input wire [23:0] pixel_data,
        input trigger,
		// Ports of Axi Master Bus Interface M00_AXIS
		input wire  m00_axis_tready,
		output logic  m00_axis_tvalid, m00_axis_tlast,
		output logic [C_M00_AXIS_TDATA_WIDTH-1 : 0] m00_axis_tdata,
		output logic [(C_M00_AXIS_TDATA_WIDTH/8)-1: 0] m00_axis_tstrb
	);
 
    //You want to send up TLAST-framed bursts of data that are 2**16 in length
    //update and test this module to make sure that's happening.
    
    logic trigger_sync[1:0];
    logic [7:0] debounce_cycles;
    logic trigger_debounced;

    logic [15:0] samples;
    logic transmitting;
    logic  handshake;
    assign handshake = transmitting && m00_axis_tready;

    always_ff @(posedge pixel_clk) begin
        trigger_sync[0] <= trigger;
        trigger_sync[1] <= trigger_sync[0]; // sync trigger and debounce below
        debounce_cycles <= (!trigger_sync[1]) ? 8'h0 : 
                           (&debounce_cycles) ? 8'b0 : debounce_cycles + 1;
        trigger_debounced       <= debounce_cycles+1'b1==8'hFF;

        transmitting <= (!transmitting && trigger_debounced) || (transmitting && !(handshake&&samples==16'hFFFF));
        samples <= (!transmitting) ? 0 : (!handshake) ? samples : (samples==16'hFFFF) ? 0 : samples + 1;
    end

    always_ff @(posedge pixel_clk) begin
        m00_axis_tvalid <= transmitting && !(samples==16'hFFFF); //?? How often should data be valid (CHANGE ME)?
        m00_axis_tlast <= handshake && samples==16'hFFFF; //when should TLAST be high (CHANGE ME)?
        m00_axis_tdata <= {8'b0, pixel_data}; //i'll give this one to you
        m00_axis_tstrb <= 4'b1111; //let's just say all bits are good all the time
    end

endmodule